module uPLogoRom (
    input logic [7:0] charAddr,
    input logic [2:0] xOffset,
    yOffset,
    output logic pixel
);
  // logic [5:0] 
endmodule
